parameter MEM_DEPTH = ;
parameter LINE_COUNT = ;